///////////////////////////////////////////////////////////////////////////////
// File:        cfs_algn_md_test_ctrlsize1_rxsize2_offset0.sv
// Author:      Pranav
// Date:        2025-07-15
// Description: Test to configure ctrl_size=1 and send RX packet with size=2, offset=0
///////////////////////////////////////////////////////////////////////////////

`ifndef CFS_ALGN_MD_TEST_CTRLSIZE1_RXSIZE2_OFFSET0_SV
`define CFS_ALGN_MD_TEST_CTRLSIZE1_RXSIZE2_OFFSET0_SV

class cfs_algn_md_test_ctrlsize1_rxsize2_offset0 extends cfs_algn_test_base;

  `uvm_component_utils(cfs_algn_md_test_ctrlsize1_rxsize2_offset0)

  function new(string name = "", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual task run_phase(uvm_phase phase);

    cfs_md_sequence_slave_response_forever resp_seq;
    cfs_algn_virtual_sequence_reg_config cfg_seq;
    cfs_algn_virtual_sequence_rx_size2_offset0 rx_seq;
    cfs_algn_virtual_sequence_rx_crt rx_seq1;
    cfs_algn_virtual_sequence_rx_size1_offset0 rx_seq2;
    cfs_algn_vif vif;
    uvm_status_e status;
    uvm_reg_data_t ctrl_val;

    phase.raise_objection(this, "TEST_START");

    #(100ns);

    // Step 0: Start slave response to keep design alive
    fork
      begin
        resp_seq = cfs_md_sequence_slave_response_forever::type_id::create("resp_seq");
        resp_seq.start(env.md_tx_agent.sequencer);
      end
    join_none

    // Step 1: Register configuration
    cfg_seq = cfs_algn_virtual_sequence_reg_config::type_id::create("cfg_seq");
    cfg_seq.set_sequencer(env.virtual_sequencer);
    cfg_seq.start(env.virtual_sequencer);

    // Step 2: Manually set CTRL: ctrl_size = 4, ctrl_offset = 0
    env.model.reg_block.CTRL.write(status, 32'h00000004, UVM_FRONTDOOR);
    env.model.reg_block.CTRL.read(status, ctrl_val, UVM_FRONTDOOR);
    `uvm_info("rxsize2_ctrlsize4", $sformatf("CTRL register value: 0x%0h", ctrl_val), UVM_MEDIUM)

    rx_seq1 = cfs_algn_virtual_sequence_rx_crt::type_id::create("rx_seq");
    rx_seq1.set_sequencer(env.virtual_sequencer);
    void'(rx_seq1.randomize());
    rx_seq1.start(env.virtual_sequencer);

    // Step 3: Send RX packet with size = 2, offset = 0 (less than ctrl_size)

    rx_seq2 = cfs_algn_virtual_sequence_rx_size1_offset0::type_id::create("rx_seq");
    rx_seq2.set_sequencer(env.virtual_sequencer);
    void'(rx_seq2.randomize());
    rx_seq2.start(env.virtual_sequencer);
    repeat (2) begin
      rx_seq = cfs_algn_virtual_sequence_rx_size2_offset0::type_id::create("rx_seq");
      rx_seq.set_sequencer(env.virtual_sequencer);
      void'(rx_seq.randomize());
      rx_seq.start(env.virtual_sequencer);
    end

    // Step 4: Wait to allow design to process

    vif = env.env_config.get_vif();

    repeat (20) @(posedge vif.clk);

    #(200ns);

    phase.drop_objection(this, "TEST_DONE");

  endtask

endclass

`endif
