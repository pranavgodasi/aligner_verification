///////////////////////////////////////////////////////////////////////////////
// File:        cfs_algn_types.sv
// Author:      Cristian Florin Slav
// Date:        2024-09-30
// Description: File  containing types required in the Aligner environment.
///////////////////////////////////////////////////////////////////////////////

`ifndef CFS_ALGN_TYPES_SV
`define CFS_ALGN_TYPES_SV

//Virtual interface
typedef virtual cfs_algn_if cfs_algn_vif;

`endif
